`default_nettype none
`timescale 1ns/1ps
module vga (
    input wire              clk
    );

endmodule

